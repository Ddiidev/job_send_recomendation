module models

@[params]
pub struct RequestText {
pub:
	to   string
	text string
}
