module types

pub type ThumbLink = string
