module services

const const_url = 'https://us.api-wa.me'
