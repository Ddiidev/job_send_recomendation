module models

@[params]
pub struct RequestImage {
pub:
	to      string
	url     string
	caption string
}
